.title KiCad schematic
.include "BC546.lib"
V1 vdd GND 5
R7 out GND 1Meg
R6 Net-_C4-Pad1_ GND 2.2k
C4 Net-_C4-Pad1_ GND 10u
Q1 Net-_C1-Pad1_ Net-_C3-Pad2_ Net-_C4-Pad1_ BC546B
R5 vdd Net-_C1-Pad1_ 2.7k
C5 Net-_C1-Pad1_ out 1u
R2 Net-_C2-Pad2_ GND 6.8k
R1 Net-_C1-Pad2_ GND 6.8k
C3 Net-_C2-Pad2_ Net-_C3-Pad2_ 2.4n
R4 Net-_C3-Pad2_ GND 6.8k
C1 Net-_C1-Pad1_ Net-_C1-Pad2_ 2.4n
C2 Net-_C1-Pad2_ Net-_C2-Pad2_ 2.4n
R3 vdd Net-_C3-Pad2_ 8.5k
.tran 10u 25m 5m
.end
