* another state machine example
* by Holger Vogt, July 9th, 2020
* 3-bit counter in a subcircuit with analog in and out

* clock
vclk cl 0 dc 0 pulse (0 5 1u 1u 1u 10u 24u)
* up or down
vupd ud 0 dc 0 pulse (0 5 1u 1u 1u 500u 1m)
* the call to the subcircuit
Xcount ud cl ob2 ob1 ob0 3bcounter


*** counter
.subckt 3bcounter updown clock out_b2 out_b1 out_b0
* Define a simple 3 bit up/down counter that counts clk edges.
* Digital outputs are on b2 b1 b0.
*   inputs  clock   reset     outputs (all digital)
a0  [upd]  clk    n_zero   [b2 b1 b0]   state2

.model state2 d_state(state_file = "state-3bit-count.in")

* Digital "one" and "zero"
a1 n_one pullup1
.model pullup1 d_pullup(load = 1pF)
a2 n_zero pulldown1
.model pulldown1 d_pulldown(load = 1pF)

* Convert the digital outputs to analog
a3 [b2] [out_b2] dac1
a4 [b1] [out_b1] dac1
a5 [b0] [out_b0] dac1
.model dac1 dac_bridge(out_low = 0 out_high = 5 out_undef = 2.5)
* Convert the analog inputs to digital
a6 [clock] [clk] adc1
a7 [updown] [upd] adc1
.model adc1 adc_bridge(in_low = 0.3 in_high = 3.5)
.ends
*** end counter

.control
tran 1us 2ms
set xbrushwidth=2
set color0=white
plot cl-12 ud-6  ob0+2*ob1+4*ob2
.endc

.end
